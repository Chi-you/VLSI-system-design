`include "./DFF.v"
`include "./4bit_cla.v"
`timescale 1ns/10ps

module Syncounter();




endmodule