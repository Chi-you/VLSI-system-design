`timescale 1ns/10ps
`include "./counter.v"

module testbench();

reg 
wire



endmodule