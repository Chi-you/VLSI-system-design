`timescale 1ns/10ps
module Counter();

input mode
output 